library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity char_rom is
	port(
		clk: in std_logic;
		char: in std_logic_vector(3 downto 0); --16 chars
		posX: in std_logic_vector(4 downto 0); -- position within the char (32x32)
		posY: in std_logic_vector(4 downto 0); -- position within the char (32x32)
		valueout: out std_logic
	);
end;

architecture behavioral of char_rom is
type rom_type is array(0 to 511) of std_logic_vector(0 to 31);
signal ROM: rom_type:= (
 0 => "00001111111111111111111100000000",	 1 => "00011111111111111111111110000000",	 2 => "00111111111111111111111111000000",	 3 => "01111111111111111111111111100000",	 4 => "11111110000000000000111111110000",	 5 => "11111100000000000001111111110000",	 6 => "11111000000000000011111111110000",	 7 => "11110000000000000111111111110000",	 8 => "11110000000000001111111011110000",	 9 => "11110000000000011111110011110000",	10 => "11110000000000111111100011110000",	11 => "11110000000001111111000011110000",	12 => "11110000000011111110000011110000",	13 => "11110000000111111100000011110000",	14 => "11110000001111111000000011110000",	15 => "11110000011111110000000011110000",	16 => "11110000111111100000000011110000",	17 => "11110001111111000000000011110000",	18 => "11110011111110000000000011110000",	19 => "11110111111100000000000011110000",	20 => "11111111111000000000000011110000",	21 => "11111111110000000000000111110000",	22 => "11111111100000000000001111110000",	23 => "11111111000000000000011111110000",	24 => "01111111111111111111111111100000",	25 => "00111111111111111111111111000000",	26 => "00011111111111111111111110000000",	27 => "00001111111111111111111100000000",	28 => "00000000000000000000000000000000",	29 => "00000000000000000000000000000000",	30 => "00000000000000000000000000000000",	31 => "00000000000000000000000000000000",	
32 => "00000000000011111000000000000000",	33 => "00000000001111111000000000000000",	34 => "00000000111111111000000000000000",	35 => "00000011111111111000000000000000",	36 => "00001111111111111000000000000000",	37 => "00001111110011111000000000000000",	38 => "00001111000011111000000000000000",	39 => "00001100000011111000000000000000",	40 => "00000000000011111000000000000000",	41 => "00000000000011111000000000000000",	42 => "00000000000011111000000000000000",	43 => "00000000000011111000000000000000",	44 => "00000000000011111000000000000000",	45 => "00000000000011111000000000000000",	46 => "00000000000011111000000000000000",	47 => "00000000000011111000000000000000",	48 => "00000000000011111000000000000000",	49 => "00000000000011111000000000000000",	50 => "00000000000011111000000000000000",	51 => "00000000000011111000000000000000",	52 => "00000000000011111000000000000000",	53 => "00000000000011111000000000000000",	54 => "00000000000011111000000000000000",	55 => "00000000000011111000000000000000",	56 => "00001111111111111111111100000000",	57 => "00001111111111111111111100000000",	58 => "00001111111111111111111100000000",	59 => "00001111111111111111111100000000",	60 => "00000000000000000000000000000000",	61 => "00000000000000000000000000000000",	62 => "00000000000000000000000000000000",	63 => "00000000000000000000000000000000",	
64 => "11111111111111111111111100000000",	65 => "11111111111111111111111110000000",	66 => "11111111111111111111111111000000",	67 => "11111111111111111111111111100000",	68 => "00000000000000000000011111110000",	69 => "00000000000000000000001111110000",	70 => "00000000000000000000000111110000",	71 => "00000000000000000000000011110000",	72 => "00000000000000000000000011110000",	73 => "00000000000000000000000011110000",	74 => "00000000000000000000000011110000",	75 => "00000000000000000000000011110000",	76 => "00001111111111111111111111110000",	77 => "00011111111111111111111111110000",	78 => "00111111111111111111111111110000",	79 => "01111111111111111111111111110000",	80 => "11111110000000000000000000000000",	81 => "11111100000000000000000000000000",	82 => "11111000000000000000000000000000",	83 => "11110000000000000000000000000000",	84 => "11110000000000000000000000000000",	85 => "11110000000000000000000000000000",	86 => "11110000000000000000000000000000",	87 => "11110000000000000000000000000000",	88 => "11111111111111111111111111110000",	89 => "11111111111111111111111111110000",	90 => "11111111111111111111111111110000",	91 => "11111111111111111111111111110000",	92 => "00000000000000000000000000000000",	93 => "00000000000000000000000000000000",	94 => "00000000000000000000000000000000",	95 => "00000000000000000000000000000000",	
96 => "11111111111111111111111100000000",	97 => "11111111111111111111111110000000",	98 => "11111111111111111111111111000000",	99 => "11111111111111111111111111100000",	100 => "00000000000000000000001111110000",	101 => "00000000000000000000000111110000",	102 => "00000000000000000000000011110000",	103 => "00000000000000000000000011110000",	104 => "00000000000000000000000011110000",	105 => "00000000000000000000000011110000",	106 => "00000000000000000000000111110000",	107 => "00000000000000000000001111110000",	108 => "11111111111111111111111111100000",	109 => "11111111111111111111111111000000",	110 => "11111111111111111111111111000000",	111 => "11111111111111111111111111100000",	112 => "00000000000000000000001111110000",	113 => "00000000000000000000000111110000",	114 => "00000000000000000000000011110000",	115 => "00000000000000000000000011110000",	116 => "00000000000000000000000011110000",	117 => "00000000000000000000000011110000",	118 => "00000000000000000000000111110000",	119 => "00000000000000000000001111110000",	120 => "11111111111111111111111111100000",	121 => "11111111111111111111111111000000",	122 => "11111111111111111111111110000000",	123 => "11111111111111111111111100000000",	124 => "00000000000000000000000000000000",	125 => "00000000000000000000000000000000",	126 => "00000000000000000000000000000000",	127 => "00000000000000000000000000000000",	
128 => "11110000000000000000000011110000",	129 => "11110000000000000000000011110000",	130 => "11110000000000000000000011110000",	131 => "11110000000000000000000011110000",	132 => "11110000000000000000000011110000",	133 => "11110000000000000000000011110000",	134 => "11110000000000000000000011110000",	135 => "11110000000000000000000011110000",	136 => "11110000000000000000000011110000",	137 => "11110000000000000000000011110000",	138 => "11111000000000000000000011110000",	139 => "11111100000000000000000011110000",	140 => "01111111111111111111111111110000",	141 => "00111111111111111111111111110000",	142 => "00011111111111111111111111110000",	143 => "00001111111111111111111111110000",	144 => "00000000000000000000000011110000",	145 => "00000000000000000000000011110000",	146 => "00000000000000000000000011110000",	147 => "00000000000000000000000011110000",	148 => "00000000000000000000000011110000",	149 => "00000000000000000000000011110000",	150 => "00000000000000000000000011110000",	151 => "00000000000000000000000011110000",	152 => "00000000000000000000000011110000",	153 => "00000000000000000000000011110000",	154 => "00000000000000000000000011110000",	155 => "00000000000000000000000011110000",	156 => "00000000000000000000000000000000",	157 => "00000000000000000000000000000000",	158 => "00000000000000000000000000000000",	159 => "00000000000000000000000000000000",	
160 => "11111111111111111111111111110000",	161 => "11111111111111111111111111110000",	162 => "11111111111111111111111111110000",	163 => "11111111111111111111111111110000",	164 => "11110000000000000000000000000000",	165 => "11110000000000000000000000000000",	166 => "11110000000000000000000000000000",	167 => "11110000000000000000000000000000",	168 => "11110000000000000000000000000000",	169 => "11110000000000000000000000000000",	170 => "11111000000000000000000000000000",	171 => "11111100000000000000000000000000",	172 => "01111111111111111111111100000000",	173 => "00111111111111111111111110000000",	174 => "00011111111111111111111111000000",	175 => "00001111111111111111111111100000",	176 => "00000000000000000000011111100000",	177 => "00000000000000000000001111100000",	178 => "00000000000000000000000111100000",	179 => "00000000000000000000000111100000",	180 => "00000000000000000000000111100000",	181 => "00000000000000000000000111100000",	182 => "00000000000000000000001111100000",	183 => "00000000000000000000011111100000",	184 => "11111111111111111111111111100000",	185 => "11111111111111111111111111000000",	186 => "11111111111111111111111110000000",	187 => "11111111111111111111111100000000",	188 => "00000000000000000000000000000000",	189 => "00000000000000000000000000000000",	190 => "00000000000000000000000000000000",	191 => "00000000000000000000000000000000",	
192 => "00001111111111111111111111110000",	193 => "00011111111111111111111111110000",	194 => "00111111111111111111111111110000",	195 => "01111111111111111111111111110000",	196 => "11111100000000000000000000000000",	197 => "11111000000000000000000000000000",	198 => "11110000000000000000000000000000",	199 => "11110000000000000000000000000000",	200 => "11110000000000000000000000000000",	201 => "11110000000000000000000000000000",	202 => "11110000000000000000000000000000",	203 => "11110000000000000000000000000000",	204 => "11111111111111111111111111000000",	205 => "11111111111111111111111111100000",	206 => "11111111111111111111111111110000",	207 => "11111111111111111111111111110000",	208 => "11110000000000000000001111110000",	209 => "11110000000000000000000111110000",	210 => "11110000000000000000000011110000",	211 => "11110000000000000000000011110000",	212 => "11110000000000000000000011110000",	213 => "11110000000000000000000011110000",	214 => "11111000000000000000000111110000",	215 => "11111100000000000000001111110000",	216 => "01111111111111111111111111100000",	217 => "00111111111111111111111111000000",	218 => "00011111111111111111111110000000",	219 => "00001111111111111111111100000000",	220 => "00000000000000000000000000000000",	221 => "00000000000000000000000000000000",	222 => "00000000000000000000000000000000",	223 => "00000000000000000000000000000000",	
224 => "00000111111111111111111111000000",	225 => "00001111111111111111111111100000",	226 => "00011111111111111111111111100000",	227 => "00111111111111111111111111100000",	228 => "00000000000000000000011111000000",	229 => "00000000000000000000011111000000",	230 => "00000000000000000000111110000000",	231 => "00000000000000000000111110000000",	232 => "00000000000000000001111100000000",	233 => "00000000000000000001111100000000",	234 => "00000000000000000011111000000000",	235 => "00000000000000000011111000000000",	236 => "00000000000000000111110000000000",	237 => "00000000000000000111110000000000",	238 => "00000000000000001111100000000000",	239 => "00000000000000001111100000000000",	240 => "00000000000000011111000000000000",	241 => "00000000000000011111000000000000",	242 => "00000000000000111110000000000000",	243 => "00000000000000111110000000000000",	244 => "00000000000001111100000000000000",	245 => "00000000000001111100000000000000",	246 => "00000000000011111000000000000000",	247 => "00000000000011111000000000000000",	248 => "00000000000111110000000000000000",	249 => "00000000000111110000000000000000",	250 => "00000000000000000000000000000000",	251 => "00000000000000000000000000000000",	252 => "00000000000000000000000000000000",	253 => "00000000000000000000000000000000",	254 => "00000000000000000000000000000000",	255 => "00000000000000000000000000000000",	
256 => "00001111111111111111111100000000",	257 => "00011111111111111111111110000000",	258 => "00111111111111111111111111000000",	259 => "01111111111111111111111111100000",	260 => "11111000000000000000000111110000",	261 => "11110000000000000000000011110000",	262 => "11110000000000000000000011110000",	263 => "11110000000000000000000011110000",	264 => "11110000000000000000000011110000",	265 => "11110000000000000000000011110000",	266 => "11110000000000000000000011110000",	267 => "11111000000000000000000111110000",	268 => "01111111111111111111111111000000",	269 => "00111111111111111111111110000000",	270 => "00111111111111111111111110000000",	271 => "01111111111111111111111111000000",	272 => "11111000000000000000000111110000",	273 => "11110000000000000000000011110000",	274 => "11110000000000000000000011110000",	275 => "11110000000000000000000011110000",	276 => "11110000000000000000000011110000",	277 => "11110000000000000000000011110000",	278 => "11110000000000000000000011110000",	279 => "11111000000000000000000111110000",	280 => "01111111111111111111111111100000",	281 => "00111111111111111111111111000000",	282 => "00011111111111111111111110000000",	283 => "00001111111111111111111100000000",	284 => "00000000000000000000000000000000",	285 => "00000000000000000000000000000000",	286 => "00000000000000000000000000000000",	287 => "00000000000000000000000000000000",	
288 => "00001111111111111111111100000000",	289 => "00011111111111111111111110000000",	290 => "00111111111111111111111111000000",	291 => "01111111111111111111111111100000",	292 => "11111100000000000000001111110000",	293 => "11111000000000000000000111110000",	294 => "11110000000000000000000011110000",	295 => "11110000000000000000000011110000",	296 => "11110000000000000000000011110000",	297 => "11110000000000000000000011110000",	298 => "11111000000000000000000011110000",	299 => "11111100000000000000000011110000",	300 => "01111111111111111111111111110000",	301 => "00111111111111111111111111110000",	302 => "00011111111111111111111111110000",	303 => "00001111111111111111111111110000",	304 => "00000000000000000000000011110000",	305 => "00000000000000000000000011110000",	306 => "00000000000000000000000011110000",	307 => "00000000000000000000000011110000",	308 => "00000000000000000000000011110000",	309 => "00000000000000000000000011110000",	310 => "00000000000000000000000111110000",	311 => "00000000000000000000001111110000",	312 => "11111111111111111111111111100000",	313 => "11111111111111111111111111000000",	314 => "11111111111111111111111110000000",	315 => "11111111111111111111111100000000",	316 => "00000000000000000000000000000000",	317 => "00000000000000000000000000000000",	318 => "00000000000000000000000000000000",	319 => "00000000000000000000000000000000",	
320 => "11110000000000000000000011110000",	321 => "11110000000000000000000011110000",	322 => "11110000000000000000000011110000",	323 => "11110000000000000000000011110000",	324 => "11110000000000000000000011110000",	325 => "11110000000000000000000011110000",	326 => "11110000000000000000000011110000",	327 => "11110000000000000000000011110000",	328 => "11110000000000000000000011110000",	329 => "11110000000000000000000011110000",	330 => "11110000000000000000000011110000",	331 => "11110000000000000000000011110000",	332 => "11110000000000000000000011110000",	333 => "11111000000000000000000111110000",	334 => "11111100000000000000001111110000",	335 => "11111110000000000000011111110000",	336 => "01111111000000000000111111100000",	337 => "00111111100000000001111111000000",	338 => "00011111110000000011111110000000",	339 => "00001111111000000111111100000000",	340 => "00000111111100001111111000000000",	341 => "00000011111110011111110000000000",	342 => "00000001111111111111100000000000",	343 => "00000000111111111111000000000000",	344 => "00000000011111111110000000000000",	345 => "00000000001111111100000000000000",	346 => "00000000000111111000000000000000",	347 => "00000000000011110000000000000000",	348 => "00000000000000000000000000000000",	349 => "00000000000000000000000000000000",	350 => "00000000000000000000000000000000",	351 => "00000000000000000000000000000000",	
352 => "00000000000000000000000000000000",	353 => "00000000000000000000000000000000",	354 => "00000000000000000000000000000000",	355 => "00000000000000000000000000000000",	356 => "00000000000000000000000000000000",	357 => "00000000000000000000000000000000",	358 => "00000000000000000000000000000000",	359 => "00000000000000000000000000000000",	360 => "00000000000000000000000000000000",	361 => "00000000000000000000000000000000",	362 => "00000000000000000000000000000000",	363 => "00000000000000000000000000000000",	364 => "00000000000000000000000000000000",	365 => "00000000000000000000000000000000",	366 => "00000000000000000000000000000000",	367 => "00000000000000000000000000000000",	368 => "00000000000011110000000000000000",	369 => "00000000000011110000000000000000",	370 => "00000000000011110000000000000000",	371 => "00000000000011110000000000000000",	372 => "00000000000011110000000000000000",	373 => "00000000000111110000000000000000",	374 => "00000000001111110000000000000000",	375 => "00000000011111110000000000000000",	376 => "00000000111111100000000000000000",	377 => "00000000111111000000000000000000",	378 => "00000000111110000000000000000000",	379 => "00000000111100000000000000000000",	380 => "00000000000000000000000000000000",	381 => "00000000000000000000000000000000",	382 => "00000000000000000000000000000000",	383 => "00000000000000000000000000000000",	
384 => "00000000000000000000000000000000",	385 => "00000000000000000000000000000000",	386 => "00000000000000000000000000000000",	387 => "00000000000000000000000000000000",	388 => "00000000000000000000000000000000",	389 => "01111000000000000010000000000000",	390 => "10000000000000000010000000000000",	391 => "10000011111001110010001110000000",	392 => "10110000010000001010010001000000",	393 => "10001000100001111010010001000000",	394 => "10001001000010001010010001000000",	395 => "01110011111001111001001110000000",	396 => "00000000000000000000000000000000",	397 => "00000000000000000000000000000000",	398 => "11110001110011110011110000000000",	399 => "00001010001000001000001000000000",	400 => "00001010011000001000001000000000",	401 => "00110010101000110011110000000000",	402 => "01000011001001000000001000000000",	403 => "10000010001010000000001000000000",	404 => "11111001110011111011110000000000",	405 => "00000000000000000000000000000000",	406 => "00000000000000000000000000000000",	407 => "00000000000000000000000000000000",	408 => "00000000000000000000000000000000",	409 => "00000000000000000000000000000000",	410 => "00000000000000000000000000000000",	411 => "00000000000000000000000000000000",	412 => "00000000000000000000000000000000",	413 => "00000000000000000000000000000000",	414 => "00000000000000000000000000000000",	415 => "00000000000000000000000000000000",	
416 => "00000000000000000000111110000000",	417 => "00000011111000000000001111111111",	418 => "00011111111001110000011111111111",	419 => "00111111111001100010011100000111",	420 => "00111110000011000010011100000111",	421 => "11100000000011000110011000000110",	422 => "11000000000110000110111000011110",	423 => "11000000000110001110110011111101",	424 => "11000000000110011110110011111101",	425 => "11000000000110111110111111100001",	426 => "11000000000111111101111111100001",	427 => "11000000000111111101100111100001",	428 => "11000000000111111101100111000001",	429 => "11000000000000011101100011000001",	430 => "11100000000000011001111111000111",	431 => "00111111100001111001111110000110",	432 => "00011111100001111001111110000110",	433 => "00000000000011100000111000001110",	434 => "00001111111111100000000000001111",	435 => "00001111111110000000000000001111",	436 => "00001111111110000000000000001111",	437 => "00000001110000000000000000000000",	438 => "00000000000000000000000000000000",	439 => "00000000000000000000000000000000",	440 => "11111110110111111101100110000110",	441 => "11111110110111111101100110000110",	442 => "11000000110111111101100110000110",	443 => "11000000110111111101100110000110",	444 => "11000000110111111101100110000110",	445 => "11000000110110011001100110000110",	446 => "11111110110110011001111110111110",	447 => "11111110110110011001111110111110",	
448 => "00000000000111111000000000000000",	449 => "00011111000110011100000000000000",	450 => "01111111000100011100000000000000",	451 => "01111000000100011100000000000000",	452 => "01110000001000011100000000000000",	453 => "01110000001001111100000000000000",	454 => "11000000111111110000000000000000",	455 => "11000000111111100000000000000000",	456 => "11000000111110000000000000000000",	457 => "10000001111110000000000000000000",	458 => "11000001111111100000000000000000",	459 => "11111001110111100000000000000000",	460 => "11111001110011100000000000000000",	461 => "00000001000001110000000000000000",	462 => "00000111000000011100000000000000",	463 => "00000111000000011110000000010000",	464 => "00000111000000001110000000010000",	465 => "00000110000000001111100000110000",	466 => "11001110000000000001111000100000",	467 => "11001110000000000001111000100000",	468 => "11001110000000000000111100100000",	469 => "00001110000000000000011111100000",	470 => "00011100000000000000000111100000",	471 => "00011100000000000000000011100000",	472 => "11111110111111111111000000100000",	473 => "11111110111100000000000000000000",	474 => "11111110111100000000000000000000",	475 => "11111110111100000000000000000000",	476 => "11111110000111110000000000000000",	477 => "11000110000111110000000000000000",	478 => "11000110111111111000000000000000",	479 => "11000110111111111000000000000000",	
480 => "00000000000000000000000000000000",	481 => "00000000000000000000000000000000",	482 => "00000000000000000000000000000000",	483 => "00000000000000000000000000000000",	484 => "00000000000000000000000000000000",	485 => "00000000000000000000000000000000",	486 => "00000000000000000000000000000000",	487 => "00000000000000000000000000000000",	488 => "00000000000000000000000000000000",	489 => "00000000000000000000000000000000",	490 => "00000000000000000000000000000000",	491 => "00000000000000000000000000000000",	492 => "00000000000000000000000000000000",	493 => "00000000000000000000000000000000",	494 => "00000000000000000000000000000000",	495 => "00000000000000000000000000000000",	496 => "00000000000000000000000000000000",	497 => "00000000000000000000000000000000",	498 => "00000000000000000000000000000000",	499 => "00000000000000000000000000000000",	500 => "00000000000000000000000000000000",	501 => "00000000000000000000000000000000",	502 => "00000000000000000000000000000000",	503 => "00000000000000000000000000000000",	504 => "00000000000000000000000000000000",	505 => "00000000000000000000000000000000",	506 => "00000000000000000000000000000000",	507 => "00000000000000000000000000000000",	508 => "00000000000000000000000000000000",	509 => "00000000000000000000000000000000",	510 => "00000000000000000000000000000000",	511 => "00000000000000000000000000000000");

signal memvalue: std_logic_vector(0 to 31);
begin
	
	process(clk)
		
	begin		
		if rising_edge(clk) then
			memvalue <= ROM(conv_integer(char & posY));
		end if;
	end process;
	
	valueout <= memvalue(conv_integer(posX));
end;